entit