library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fpga_top is
port (
    -- --------------------------------
    -- CLOCKS
    ----------------------------------- 
    -- Reference clocks
    CLK		: in std_logic;
    -- Reset button
    RESET   : in std_logic; 
    
    -- --------------------------------
    -- UART
    -- --------------------------------
    -- TODO
);
end entity;

architecture full of fpga_top is
	signal clk_c0 		: std_logic;
	signal reset_cnt	: unsigned(6 downto 0);
    signal locked		: std_logic;
    signal reset_c0 	: std_logic	:= '1';

    signal btn_debounced_n      : std_logic;
    signal btn_debounced        : std_logic;
	
begin

    -- ------------------------------------------------------------------------
    -- Clocks & Reset
    -- ------------------------------------------------------------------------

    -- Clocks are generated by the PLL from reference closk 12MHz. The reset is
    -- asserted automatically when the output clocks are locked. There is also a 
    -- possibility to assert the system reset by the reset buttton.
    --
    -- List of generated clocks & resets:
    -- * clk_c0 and reset_c0 -- main system clocks used in the design

    -- Generate input clocks
    pll_i : work.pll 
    port map(
        inclk0		=> CLK,
        c0			=> clk_c0,
        locked		=> locked
    );

    -- Debounce the reset button 
    debounce_i : work.debounce
    generic map (
        counter_size  => 19
    )
    port map (
        clk     => clk_c0,
        button  => BTN,
        result  => btn_debounced_n
    );

    -- Output value from the debouncer is inverted
    btn_debounced <= not(btn_debounced_n);

    -- Reset generation is based on the counter which holds the reset for 
    -- several clock cycles. The generator of the funciton is taken from the
    -- MSB bit of the counter vector.
    reset_p : process(clk_c0)
    begin
        if(rising_edge(clk_c0))then
            if(locked = '0' or btn_debounced = '0') then
                -- Reset is locked
                reset_cnt  <= (others=>'0');
            else
                -- Reset needs to be asserted (one clock cycle shoudl be enough)
                if(reset_cnt(6) = '0')then
                    reset_cnt <= reset_cnt + 1;
                end if;
            end if;
        end if;
    end process;

    -- Output reset signal
    reset_c0 <= not(reset_cnt(6));

    -- ------------------------------------------------------------------------
    -- UART connection
    -- ------------------------------------------------------------------------
	
end architecture;
